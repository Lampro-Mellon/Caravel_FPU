magic
tech sky130A
magscale 1 2
timestamp 1623744702
<< obsli1 >>
rect 1104 17 178848 117521
<< obsm1 >>
rect 106 8 179846 117552
<< metal2 >>
rect 754 119200 810 120000
rect 2318 119200 2374 120000
rect 3882 119200 3938 120000
rect 5446 119200 5502 120000
rect 7010 119200 7066 120000
rect 8574 119200 8630 120000
rect 10138 119200 10194 120000
rect 11702 119200 11758 120000
rect 13266 119200 13322 120000
rect 14830 119200 14886 120000
rect 16394 119200 16450 120000
rect 17958 119200 18014 120000
rect 19522 119200 19578 120000
rect 21086 119200 21142 120000
rect 22650 119200 22706 120000
rect 24214 119200 24270 120000
rect 25778 119200 25834 120000
rect 27342 119200 27398 120000
rect 28906 119200 28962 120000
rect 30470 119200 30526 120000
rect 32034 119200 32090 120000
rect 33598 119200 33654 120000
rect 35162 119200 35218 120000
rect 36726 119200 36782 120000
rect 38290 119200 38346 120000
rect 39854 119200 39910 120000
rect 41418 119200 41474 120000
rect 42982 119200 43038 120000
rect 44546 119200 44602 120000
rect 46110 119200 46166 120000
rect 47674 119200 47730 120000
rect 49238 119200 49294 120000
rect 50802 119200 50858 120000
rect 52366 119200 52422 120000
rect 53930 119200 53986 120000
rect 55494 119200 55550 120000
rect 57058 119200 57114 120000
rect 58622 119200 58678 120000
rect 60186 119200 60242 120000
rect 61750 119200 61806 120000
rect 63314 119200 63370 120000
rect 64878 119200 64934 120000
rect 66442 119200 66498 120000
rect 68006 119200 68062 120000
rect 69570 119200 69626 120000
rect 71134 119200 71190 120000
rect 72698 119200 72754 120000
rect 74262 119200 74318 120000
rect 75826 119200 75882 120000
rect 77390 119200 77446 120000
rect 78954 119200 79010 120000
rect 80518 119200 80574 120000
rect 82082 119200 82138 120000
rect 83646 119200 83702 120000
rect 85210 119200 85266 120000
rect 86774 119200 86830 120000
rect 88338 119200 88394 120000
rect 89902 119200 89958 120000
rect 91558 119200 91614 120000
rect 93122 119200 93178 120000
rect 94686 119200 94742 120000
rect 96250 119200 96306 120000
rect 97814 119200 97870 120000
rect 99378 119200 99434 120000
rect 100942 119200 100998 120000
rect 102506 119200 102562 120000
rect 104070 119200 104126 120000
rect 105634 119200 105690 120000
rect 107198 119200 107254 120000
rect 108762 119200 108818 120000
rect 110326 119200 110382 120000
rect 111890 119200 111946 120000
rect 113454 119200 113510 120000
rect 115018 119200 115074 120000
rect 116582 119200 116638 120000
rect 118146 119200 118202 120000
rect 119710 119200 119766 120000
rect 121274 119200 121330 120000
rect 122838 119200 122894 120000
rect 124402 119200 124458 120000
rect 125966 119200 126022 120000
rect 127530 119200 127586 120000
rect 129094 119200 129150 120000
rect 130658 119200 130714 120000
rect 132222 119200 132278 120000
rect 133786 119200 133842 120000
rect 135350 119200 135406 120000
rect 136914 119200 136970 120000
rect 138478 119200 138534 120000
rect 140042 119200 140098 120000
rect 141606 119200 141662 120000
rect 143170 119200 143226 120000
rect 144734 119200 144790 120000
rect 146298 119200 146354 120000
rect 147862 119200 147918 120000
rect 149426 119200 149482 120000
rect 150990 119200 151046 120000
rect 152554 119200 152610 120000
rect 154118 119200 154174 120000
rect 155682 119200 155738 120000
rect 157246 119200 157302 120000
rect 158810 119200 158866 120000
rect 160374 119200 160430 120000
rect 161938 119200 161994 120000
rect 163502 119200 163558 120000
rect 165066 119200 165122 120000
rect 166630 119200 166686 120000
rect 168194 119200 168250 120000
rect 169758 119200 169814 120000
rect 171322 119200 171378 120000
rect 172886 119200 172942 120000
rect 174450 119200 174506 120000
rect 176014 119200 176070 120000
rect 177578 119200 177634 120000
rect 179142 119200 179198 120000
rect 110 0 166 800
rect 386 0 442 800
rect 754 0 810 800
rect 1122 0 1178 800
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 4066 0 4122 800
rect 4434 0 4490 800
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5538 0 5594 800
rect 5906 0 5962 800
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 7010 0 7066 800
rect 7378 0 7434 800
rect 7746 0 7802 800
rect 8114 0 8170 800
rect 8482 0 8538 800
rect 8850 0 8906 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 9954 0 10010 800
rect 10322 0 10378 800
rect 10690 0 10746 800
rect 11058 0 11114 800
rect 11426 0 11482 800
rect 11794 0 11850 800
rect 12162 0 12218 800
rect 12530 0 12586 800
rect 12898 0 12954 800
rect 13266 0 13322 800
rect 13634 0 13690 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15106 0 15162 800
rect 15474 0 15530 800
rect 15842 0 15898 800
rect 16210 0 16266 800
rect 16486 0 16542 800
rect 16854 0 16910 800
rect 17222 0 17278 800
rect 17590 0 17646 800
rect 17958 0 18014 800
rect 18326 0 18382 800
rect 18694 0 18750 800
rect 19062 0 19118 800
rect 19430 0 19486 800
rect 19798 0 19854 800
rect 20166 0 20222 800
rect 20534 0 20590 800
rect 20902 0 20958 800
rect 21270 0 21326 800
rect 21638 0 21694 800
rect 22006 0 22062 800
rect 22374 0 22430 800
rect 22742 0 22798 800
rect 23110 0 23166 800
rect 23478 0 23534 800
rect 23846 0 23902 800
rect 24214 0 24270 800
rect 24582 0 24638 800
rect 24950 0 25006 800
rect 25318 0 25374 800
rect 25686 0 25742 800
rect 26054 0 26110 800
rect 26422 0 26478 800
rect 26790 0 26846 800
rect 27158 0 27214 800
rect 27526 0 27582 800
rect 27894 0 27950 800
rect 28262 0 28318 800
rect 28630 0 28686 800
rect 28998 0 29054 800
rect 29366 0 29422 800
rect 29734 0 29790 800
rect 30102 0 30158 800
rect 30470 0 30526 800
rect 30838 0 30894 800
rect 31206 0 31262 800
rect 31574 0 31630 800
rect 31942 0 31998 800
rect 32310 0 32366 800
rect 32678 0 32734 800
rect 32954 0 33010 800
rect 33322 0 33378 800
rect 33690 0 33746 800
rect 34058 0 34114 800
rect 34426 0 34482 800
rect 34794 0 34850 800
rect 35162 0 35218 800
rect 35530 0 35586 800
rect 35898 0 35954 800
rect 36266 0 36322 800
rect 36634 0 36690 800
rect 37002 0 37058 800
rect 37370 0 37426 800
rect 37738 0 37794 800
rect 38106 0 38162 800
rect 38474 0 38530 800
rect 38842 0 38898 800
rect 39210 0 39266 800
rect 39578 0 39634 800
rect 39946 0 40002 800
rect 40314 0 40370 800
rect 40682 0 40738 800
rect 41050 0 41106 800
rect 41418 0 41474 800
rect 41786 0 41842 800
rect 42154 0 42210 800
rect 42522 0 42578 800
rect 42890 0 42946 800
rect 43258 0 43314 800
rect 43626 0 43682 800
rect 43994 0 44050 800
rect 44362 0 44418 800
rect 44730 0 44786 800
rect 45098 0 45154 800
rect 45466 0 45522 800
rect 45834 0 45890 800
rect 46202 0 46258 800
rect 46570 0 46626 800
rect 46938 0 46994 800
rect 47306 0 47362 800
rect 47674 0 47730 800
rect 48042 0 48098 800
rect 48410 0 48466 800
rect 48778 0 48834 800
rect 49146 0 49202 800
rect 49422 0 49478 800
rect 49790 0 49846 800
rect 50158 0 50214 800
rect 50526 0 50582 800
rect 50894 0 50950 800
rect 51262 0 51318 800
rect 51630 0 51686 800
rect 51998 0 52054 800
rect 52366 0 52422 800
rect 52734 0 52790 800
rect 53102 0 53158 800
rect 53470 0 53526 800
rect 53838 0 53894 800
rect 54206 0 54262 800
rect 54574 0 54630 800
rect 54942 0 54998 800
rect 55310 0 55366 800
rect 55678 0 55734 800
rect 56046 0 56102 800
rect 56414 0 56470 800
rect 56782 0 56838 800
rect 57150 0 57206 800
rect 57518 0 57574 800
rect 57886 0 57942 800
rect 58254 0 58310 800
rect 58622 0 58678 800
rect 58990 0 59046 800
rect 59358 0 59414 800
rect 59726 0 59782 800
rect 60094 0 60150 800
rect 60462 0 60518 800
rect 60830 0 60886 800
rect 61198 0 61254 800
rect 61566 0 61622 800
rect 61934 0 61990 800
rect 62302 0 62358 800
rect 62670 0 62726 800
rect 63038 0 63094 800
rect 63406 0 63462 800
rect 63774 0 63830 800
rect 64142 0 64198 800
rect 64510 0 64566 800
rect 64878 0 64934 800
rect 65246 0 65302 800
rect 65522 0 65578 800
rect 65890 0 65946 800
rect 66258 0 66314 800
rect 66626 0 66682 800
rect 66994 0 67050 800
rect 67362 0 67418 800
rect 67730 0 67786 800
rect 68098 0 68154 800
rect 68466 0 68522 800
rect 68834 0 68890 800
rect 69202 0 69258 800
rect 69570 0 69626 800
rect 69938 0 69994 800
rect 70306 0 70362 800
rect 70674 0 70730 800
rect 71042 0 71098 800
rect 71410 0 71466 800
rect 71778 0 71834 800
rect 72146 0 72202 800
rect 72514 0 72570 800
rect 72882 0 72938 800
rect 73250 0 73306 800
rect 73618 0 73674 800
rect 73986 0 74042 800
rect 74354 0 74410 800
rect 74722 0 74778 800
rect 75090 0 75146 800
rect 75458 0 75514 800
rect 75826 0 75882 800
rect 76194 0 76250 800
rect 76562 0 76618 800
rect 76930 0 76986 800
rect 77298 0 77354 800
rect 77666 0 77722 800
rect 78034 0 78090 800
rect 78402 0 78458 800
rect 78770 0 78826 800
rect 79138 0 79194 800
rect 79506 0 79562 800
rect 79874 0 79930 800
rect 80242 0 80298 800
rect 80610 0 80666 800
rect 80978 0 81034 800
rect 81346 0 81402 800
rect 81714 0 81770 800
rect 81990 0 82046 800
rect 82358 0 82414 800
rect 82726 0 82782 800
rect 83094 0 83150 800
rect 83462 0 83518 800
rect 83830 0 83886 800
rect 84198 0 84254 800
rect 84566 0 84622 800
rect 84934 0 84990 800
rect 85302 0 85358 800
rect 85670 0 85726 800
rect 86038 0 86094 800
rect 86406 0 86462 800
rect 86774 0 86830 800
rect 87142 0 87198 800
rect 87510 0 87566 800
rect 87878 0 87934 800
rect 88246 0 88302 800
rect 88614 0 88670 800
rect 88982 0 89038 800
rect 89350 0 89406 800
rect 89718 0 89774 800
rect 90086 0 90142 800
rect 90454 0 90510 800
rect 90822 0 90878 800
rect 91190 0 91246 800
rect 91558 0 91614 800
rect 91926 0 91982 800
rect 92294 0 92350 800
rect 92662 0 92718 800
rect 93030 0 93086 800
rect 93398 0 93454 800
rect 93766 0 93822 800
rect 94134 0 94190 800
rect 94502 0 94558 800
rect 94870 0 94926 800
rect 95238 0 95294 800
rect 95606 0 95662 800
rect 95974 0 96030 800
rect 96342 0 96398 800
rect 96710 0 96766 800
rect 97078 0 97134 800
rect 97446 0 97502 800
rect 97814 0 97870 800
rect 98182 0 98238 800
rect 98458 0 98514 800
rect 98826 0 98882 800
rect 99194 0 99250 800
rect 99562 0 99618 800
rect 99930 0 99986 800
rect 100298 0 100354 800
rect 100666 0 100722 800
rect 101034 0 101090 800
rect 101402 0 101458 800
rect 101770 0 101826 800
rect 102138 0 102194 800
rect 102506 0 102562 800
rect 102874 0 102930 800
rect 103242 0 103298 800
rect 103610 0 103666 800
rect 103978 0 104034 800
rect 104346 0 104402 800
rect 104714 0 104770 800
rect 105082 0 105138 800
rect 105450 0 105506 800
rect 105818 0 105874 800
rect 106186 0 106242 800
rect 106554 0 106610 800
rect 106922 0 106978 800
rect 107290 0 107346 800
rect 107658 0 107714 800
rect 108026 0 108082 800
rect 108394 0 108450 800
rect 108762 0 108818 800
rect 109130 0 109186 800
rect 109498 0 109554 800
rect 109866 0 109922 800
rect 110234 0 110290 800
rect 110602 0 110658 800
rect 110970 0 111026 800
rect 111338 0 111394 800
rect 111706 0 111762 800
rect 112074 0 112130 800
rect 112442 0 112498 800
rect 112810 0 112866 800
rect 113178 0 113234 800
rect 113546 0 113602 800
rect 113914 0 113970 800
rect 114282 0 114338 800
rect 114650 0 114706 800
rect 114926 0 114982 800
rect 115294 0 115350 800
rect 115662 0 115718 800
rect 116030 0 116086 800
rect 116398 0 116454 800
rect 116766 0 116822 800
rect 117134 0 117190 800
rect 117502 0 117558 800
rect 117870 0 117926 800
rect 118238 0 118294 800
rect 118606 0 118662 800
rect 118974 0 119030 800
rect 119342 0 119398 800
rect 119710 0 119766 800
rect 120078 0 120134 800
rect 120446 0 120502 800
rect 120814 0 120870 800
rect 121182 0 121238 800
rect 121550 0 121606 800
rect 121918 0 121974 800
rect 122286 0 122342 800
rect 122654 0 122710 800
rect 123022 0 123078 800
rect 123390 0 123446 800
rect 123758 0 123814 800
rect 124126 0 124182 800
rect 124494 0 124550 800
rect 124862 0 124918 800
rect 125230 0 125286 800
rect 125598 0 125654 800
rect 125966 0 126022 800
rect 126334 0 126390 800
rect 126702 0 126758 800
rect 127070 0 127126 800
rect 127438 0 127494 800
rect 127806 0 127862 800
rect 128174 0 128230 800
rect 128542 0 128598 800
rect 128910 0 128966 800
rect 129278 0 129334 800
rect 129646 0 129702 800
rect 130014 0 130070 800
rect 130382 0 130438 800
rect 130750 0 130806 800
rect 131026 0 131082 800
rect 131394 0 131450 800
rect 131762 0 131818 800
rect 132130 0 132186 800
rect 132498 0 132554 800
rect 132866 0 132922 800
rect 133234 0 133290 800
rect 133602 0 133658 800
rect 133970 0 134026 800
rect 134338 0 134394 800
rect 134706 0 134762 800
rect 135074 0 135130 800
rect 135442 0 135498 800
rect 135810 0 135866 800
rect 136178 0 136234 800
rect 136546 0 136602 800
rect 136914 0 136970 800
rect 137282 0 137338 800
rect 137650 0 137706 800
rect 138018 0 138074 800
rect 138386 0 138442 800
rect 138754 0 138810 800
rect 139122 0 139178 800
rect 139490 0 139546 800
rect 139858 0 139914 800
rect 140226 0 140282 800
rect 140594 0 140650 800
rect 140962 0 141018 800
rect 141330 0 141386 800
rect 141698 0 141754 800
rect 142066 0 142122 800
rect 142434 0 142490 800
rect 142802 0 142858 800
rect 143170 0 143226 800
rect 143538 0 143594 800
rect 143906 0 143962 800
rect 144274 0 144330 800
rect 144642 0 144698 800
rect 145010 0 145066 800
rect 145378 0 145434 800
rect 145746 0 145802 800
rect 146114 0 146170 800
rect 146482 0 146538 800
rect 146850 0 146906 800
rect 147218 0 147274 800
rect 147494 0 147550 800
rect 147862 0 147918 800
rect 148230 0 148286 800
rect 148598 0 148654 800
rect 148966 0 149022 800
rect 149334 0 149390 800
rect 149702 0 149758 800
rect 150070 0 150126 800
rect 150438 0 150494 800
rect 150806 0 150862 800
rect 151174 0 151230 800
rect 151542 0 151598 800
rect 151910 0 151966 800
rect 152278 0 152334 800
rect 152646 0 152702 800
rect 153014 0 153070 800
rect 153382 0 153438 800
rect 153750 0 153806 800
rect 154118 0 154174 800
rect 154486 0 154542 800
rect 154854 0 154910 800
rect 155222 0 155278 800
rect 155590 0 155646 800
rect 155958 0 156014 800
rect 156326 0 156382 800
rect 156694 0 156750 800
rect 157062 0 157118 800
rect 157430 0 157486 800
rect 157798 0 157854 800
rect 158166 0 158222 800
rect 158534 0 158590 800
rect 158902 0 158958 800
rect 159270 0 159326 800
rect 159638 0 159694 800
rect 160006 0 160062 800
rect 160374 0 160430 800
rect 160742 0 160798 800
rect 161110 0 161166 800
rect 161478 0 161534 800
rect 161846 0 161902 800
rect 162214 0 162270 800
rect 162582 0 162638 800
rect 162950 0 163006 800
rect 163318 0 163374 800
rect 163686 0 163742 800
rect 163962 0 164018 800
rect 164330 0 164386 800
rect 164698 0 164754 800
rect 165066 0 165122 800
rect 165434 0 165490 800
rect 165802 0 165858 800
rect 166170 0 166226 800
rect 166538 0 166594 800
rect 166906 0 166962 800
rect 167274 0 167330 800
rect 167642 0 167698 800
rect 168010 0 168066 800
rect 168378 0 168434 800
rect 168746 0 168802 800
rect 169114 0 169170 800
rect 169482 0 169538 800
rect 169850 0 169906 800
rect 170218 0 170274 800
rect 170586 0 170642 800
rect 170954 0 171010 800
rect 171322 0 171378 800
rect 171690 0 171746 800
rect 172058 0 172114 800
rect 172426 0 172482 800
rect 172794 0 172850 800
rect 173162 0 173218 800
rect 173530 0 173586 800
rect 173898 0 173954 800
rect 174266 0 174322 800
rect 174634 0 174690 800
rect 175002 0 175058 800
rect 175370 0 175426 800
rect 175738 0 175794 800
rect 176106 0 176162 800
rect 176474 0 176530 800
rect 176842 0 176898 800
rect 177210 0 177266 800
rect 177578 0 177634 800
rect 177946 0 178002 800
rect 178314 0 178370 800
rect 178682 0 178738 800
rect 179050 0 179106 800
rect 179418 0 179474 800
rect 179786 0 179842 800
<< obsm2 >>
rect 112 119144 698 119200
rect 866 119144 2262 119200
rect 2430 119144 3826 119200
rect 3994 119144 5390 119200
rect 5558 119144 6954 119200
rect 7122 119144 8518 119200
rect 8686 119144 10082 119200
rect 10250 119144 11646 119200
rect 11814 119144 13210 119200
rect 13378 119144 14774 119200
rect 14942 119144 16338 119200
rect 16506 119144 17902 119200
rect 18070 119144 19466 119200
rect 19634 119144 21030 119200
rect 21198 119144 22594 119200
rect 22762 119144 24158 119200
rect 24326 119144 25722 119200
rect 25890 119144 27286 119200
rect 27454 119144 28850 119200
rect 29018 119144 30414 119200
rect 30582 119144 31978 119200
rect 32146 119144 33542 119200
rect 33710 119144 35106 119200
rect 35274 119144 36670 119200
rect 36838 119144 38234 119200
rect 38402 119144 39798 119200
rect 39966 119144 41362 119200
rect 41530 119144 42926 119200
rect 43094 119144 44490 119200
rect 44658 119144 46054 119200
rect 46222 119144 47618 119200
rect 47786 119144 49182 119200
rect 49350 119144 50746 119200
rect 50914 119144 52310 119200
rect 52478 119144 53874 119200
rect 54042 119144 55438 119200
rect 55606 119144 57002 119200
rect 57170 119144 58566 119200
rect 58734 119144 60130 119200
rect 60298 119144 61694 119200
rect 61862 119144 63258 119200
rect 63426 119144 64822 119200
rect 64990 119144 66386 119200
rect 66554 119144 67950 119200
rect 68118 119144 69514 119200
rect 69682 119144 71078 119200
rect 71246 119144 72642 119200
rect 72810 119144 74206 119200
rect 74374 119144 75770 119200
rect 75938 119144 77334 119200
rect 77502 119144 78898 119200
rect 79066 119144 80462 119200
rect 80630 119144 82026 119200
rect 82194 119144 83590 119200
rect 83758 119144 85154 119200
rect 85322 119144 86718 119200
rect 86886 119144 88282 119200
rect 88450 119144 89846 119200
rect 90014 119144 91502 119200
rect 91670 119144 93066 119200
rect 93234 119144 94630 119200
rect 94798 119144 96194 119200
rect 96362 119144 97758 119200
rect 97926 119144 99322 119200
rect 99490 119144 100886 119200
rect 101054 119144 102450 119200
rect 102618 119144 104014 119200
rect 104182 119144 105578 119200
rect 105746 119144 107142 119200
rect 107310 119144 108706 119200
rect 108874 119144 110270 119200
rect 110438 119144 111834 119200
rect 112002 119144 113398 119200
rect 113566 119144 114962 119200
rect 115130 119144 116526 119200
rect 116694 119144 118090 119200
rect 118258 119144 119654 119200
rect 119822 119144 121218 119200
rect 121386 119144 122782 119200
rect 122950 119144 124346 119200
rect 124514 119144 125910 119200
rect 126078 119144 127474 119200
rect 127642 119144 129038 119200
rect 129206 119144 130602 119200
rect 130770 119144 132166 119200
rect 132334 119144 133730 119200
rect 133898 119144 135294 119200
rect 135462 119144 136858 119200
rect 137026 119144 138422 119200
rect 138590 119144 139986 119200
rect 140154 119144 141550 119200
rect 141718 119144 143114 119200
rect 143282 119144 144678 119200
rect 144846 119144 146242 119200
rect 146410 119144 147806 119200
rect 147974 119144 149370 119200
rect 149538 119144 150934 119200
rect 151102 119144 152498 119200
rect 152666 119144 154062 119200
rect 154230 119144 155626 119200
rect 155794 119144 157190 119200
rect 157358 119144 158754 119200
rect 158922 119144 160318 119200
rect 160486 119144 161882 119200
rect 162050 119144 163446 119200
rect 163614 119144 165010 119200
rect 165178 119144 166574 119200
rect 166742 119144 168138 119200
rect 168306 119144 169702 119200
rect 169870 119144 171266 119200
rect 171434 119144 172830 119200
rect 172998 119144 174394 119200
rect 174562 119144 175958 119200
rect 176126 119144 177522 119200
rect 177690 119144 179086 119200
rect 179254 119144 179840 119200
rect 112 856 179840 119144
rect 222 2 330 856
rect 498 2 698 856
rect 866 2 1066 856
rect 1234 2 1434 856
rect 1602 2 1802 856
rect 1970 2 2170 856
rect 2338 2 2538 856
rect 2706 2 2906 856
rect 3074 2 3274 856
rect 3442 2 3642 856
rect 3810 2 4010 856
rect 4178 2 4378 856
rect 4546 2 4746 856
rect 4914 2 5114 856
rect 5282 2 5482 856
rect 5650 2 5850 856
rect 6018 2 6218 856
rect 6386 2 6586 856
rect 6754 2 6954 856
rect 7122 2 7322 856
rect 7490 2 7690 856
rect 7858 2 8058 856
rect 8226 2 8426 856
rect 8594 2 8794 856
rect 8962 2 9162 856
rect 9330 2 9530 856
rect 9698 2 9898 856
rect 10066 2 10266 856
rect 10434 2 10634 856
rect 10802 2 11002 856
rect 11170 2 11370 856
rect 11538 2 11738 856
rect 11906 2 12106 856
rect 12274 2 12474 856
rect 12642 2 12842 856
rect 13010 2 13210 856
rect 13378 2 13578 856
rect 13746 2 13946 856
rect 14114 2 14314 856
rect 14482 2 14682 856
rect 14850 2 15050 856
rect 15218 2 15418 856
rect 15586 2 15786 856
rect 15954 2 16154 856
rect 16322 2 16430 856
rect 16598 2 16798 856
rect 16966 2 17166 856
rect 17334 2 17534 856
rect 17702 2 17902 856
rect 18070 2 18270 856
rect 18438 2 18638 856
rect 18806 2 19006 856
rect 19174 2 19374 856
rect 19542 2 19742 856
rect 19910 2 20110 856
rect 20278 2 20478 856
rect 20646 2 20846 856
rect 21014 2 21214 856
rect 21382 2 21582 856
rect 21750 2 21950 856
rect 22118 2 22318 856
rect 22486 2 22686 856
rect 22854 2 23054 856
rect 23222 2 23422 856
rect 23590 2 23790 856
rect 23958 2 24158 856
rect 24326 2 24526 856
rect 24694 2 24894 856
rect 25062 2 25262 856
rect 25430 2 25630 856
rect 25798 2 25998 856
rect 26166 2 26366 856
rect 26534 2 26734 856
rect 26902 2 27102 856
rect 27270 2 27470 856
rect 27638 2 27838 856
rect 28006 2 28206 856
rect 28374 2 28574 856
rect 28742 2 28942 856
rect 29110 2 29310 856
rect 29478 2 29678 856
rect 29846 2 30046 856
rect 30214 2 30414 856
rect 30582 2 30782 856
rect 30950 2 31150 856
rect 31318 2 31518 856
rect 31686 2 31886 856
rect 32054 2 32254 856
rect 32422 2 32622 856
rect 32790 2 32898 856
rect 33066 2 33266 856
rect 33434 2 33634 856
rect 33802 2 34002 856
rect 34170 2 34370 856
rect 34538 2 34738 856
rect 34906 2 35106 856
rect 35274 2 35474 856
rect 35642 2 35842 856
rect 36010 2 36210 856
rect 36378 2 36578 856
rect 36746 2 36946 856
rect 37114 2 37314 856
rect 37482 2 37682 856
rect 37850 2 38050 856
rect 38218 2 38418 856
rect 38586 2 38786 856
rect 38954 2 39154 856
rect 39322 2 39522 856
rect 39690 2 39890 856
rect 40058 2 40258 856
rect 40426 2 40626 856
rect 40794 2 40994 856
rect 41162 2 41362 856
rect 41530 2 41730 856
rect 41898 2 42098 856
rect 42266 2 42466 856
rect 42634 2 42834 856
rect 43002 2 43202 856
rect 43370 2 43570 856
rect 43738 2 43938 856
rect 44106 2 44306 856
rect 44474 2 44674 856
rect 44842 2 45042 856
rect 45210 2 45410 856
rect 45578 2 45778 856
rect 45946 2 46146 856
rect 46314 2 46514 856
rect 46682 2 46882 856
rect 47050 2 47250 856
rect 47418 2 47618 856
rect 47786 2 47986 856
rect 48154 2 48354 856
rect 48522 2 48722 856
rect 48890 2 49090 856
rect 49258 2 49366 856
rect 49534 2 49734 856
rect 49902 2 50102 856
rect 50270 2 50470 856
rect 50638 2 50838 856
rect 51006 2 51206 856
rect 51374 2 51574 856
rect 51742 2 51942 856
rect 52110 2 52310 856
rect 52478 2 52678 856
rect 52846 2 53046 856
rect 53214 2 53414 856
rect 53582 2 53782 856
rect 53950 2 54150 856
rect 54318 2 54518 856
rect 54686 2 54886 856
rect 55054 2 55254 856
rect 55422 2 55622 856
rect 55790 2 55990 856
rect 56158 2 56358 856
rect 56526 2 56726 856
rect 56894 2 57094 856
rect 57262 2 57462 856
rect 57630 2 57830 856
rect 57998 2 58198 856
rect 58366 2 58566 856
rect 58734 2 58934 856
rect 59102 2 59302 856
rect 59470 2 59670 856
rect 59838 2 60038 856
rect 60206 2 60406 856
rect 60574 2 60774 856
rect 60942 2 61142 856
rect 61310 2 61510 856
rect 61678 2 61878 856
rect 62046 2 62246 856
rect 62414 2 62614 856
rect 62782 2 62982 856
rect 63150 2 63350 856
rect 63518 2 63718 856
rect 63886 2 64086 856
rect 64254 2 64454 856
rect 64622 2 64822 856
rect 64990 2 65190 856
rect 65358 2 65466 856
rect 65634 2 65834 856
rect 66002 2 66202 856
rect 66370 2 66570 856
rect 66738 2 66938 856
rect 67106 2 67306 856
rect 67474 2 67674 856
rect 67842 2 68042 856
rect 68210 2 68410 856
rect 68578 2 68778 856
rect 68946 2 69146 856
rect 69314 2 69514 856
rect 69682 2 69882 856
rect 70050 2 70250 856
rect 70418 2 70618 856
rect 70786 2 70986 856
rect 71154 2 71354 856
rect 71522 2 71722 856
rect 71890 2 72090 856
rect 72258 2 72458 856
rect 72626 2 72826 856
rect 72994 2 73194 856
rect 73362 2 73562 856
rect 73730 2 73930 856
rect 74098 2 74298 856
rect 74466 2 74666 856
rect 74834 2 75034 856
rect 75202 2 75402 856
rect 75570 2 75770 856
rect 75938 2 76138 856
rect 76306 2 76506 856
rect 76674 2 76874 856
rect 77042 2 77242 856
rect 77410 2 77610 856
rect 77778 2 77978 856
rect 78146 2 78346 856
rect 78514 2 78714 856
rect 78882 2 79082 856
rect 79250 2 79450 856
rect 79618 2 79818 856
rect 79986 2 80186 856
rect 80354 2 80554 856
rect 80722 2 80922 856
rect 81090 2 81290 856
rect 81458 2 81658 856
rect 81826 2 81934 856
rect 82102 2 82302 856
rect 82470 2 82670 856
rect 82838 2 83038 856
rect 83206 2 83406 856
rect 83574 2 83774 856
rect 83942 2 84142 856
rect 84310 2 84510 856
rect 84678 2 84878 856
rect 85046 2 85246 856
rect 85414 2 85614 856
rect 85782 2 85982 856
rect 86150 2 86350 856
rect 86518 2 86718 856
rect 86886 2 87086 856
rect 87254 2 87454 856
rect 87622 2 87822 856
rect 87990 2 88190 856
rect 88358 2 88558 856
rect 88726 2 88926 856
rect 89094 2 89294 856
rect 89462 2 89662 856
rect 89830 2 90030 856
rect 90198 2 90398 856
rect 90566 2 90766 856
rect 90934 2 91134 856
rect 91302 2 91502 856
rect 91670 2 91870 856
rect 92038 2 92238 856
rect 92406 2 92606 856
rect 92774 2 92974 856
rect 93142 2 93342 856
rect 93510 2 93710 856
rect 93878 2 94078 856
rect 94246 2 94446 856
rect 94614 2 94814 856
rect 94982 2 95182 856
rect 95350 2 95550 856
rect 95718 2 95918 856
rect 96086 2 96286 856
rect 96454 2 96654 856
rect 96822 2 97022 856
rect 97190 2 97390 856
rect 97558 2 97758 856
rect 97926 2 98126 856
rect 98294 2 98402 856
rect 98570 2 98770 856
rect 98938 2 99138 856
rect 99306 2 99506 856
rect 99674 2 99874 856
rect 100042 2 100242 856
rect 100410 2 100610 856
rect 100778 2 100978 856
rect 101146 2 101346 856
rect 101514 2 101714 856
rect 101882 2 102082 856
rect 102250 2 102450 856
rect 102618 2 102818 856
rect 102986 2 103186 856
rect 103354 2 103554 856
rect 103722 2 103922 856
rect 104090 2 104290 856
rect 104458 2 104658 856
rect 104826 2 105026 856
rect 105194 2 105394 856
rect 105562 2 105762 856
rect 105930 2 106130 856
rect 106298 2 106498 856
rect 106666 2 106866 856
rect 107034 2 107234 856
rect 107402 2 107602 856
rect 107770 2 107970 856
rect 108138 2 108338 856
rect 108506 2 108706 856
rect 108874 2 109074 856
rect 109242 2 109442 856
rect 109610 2 109810 856
rect 109978 2 110178 856
rect 110346 2 110546 856
rect 110714 2 110914 856
rect 111082 2 111282 856
rect 111450 2 111650 856
rect 111818 2 112018 856
rect 112186 2 112386 856
rect 112554 2 112754 856
rect 112922 2 113122 856
rect 113290 2 113490 856
rect 113658 2 113858 856
rect 114026 2 114226 856
rect 114394 2 114594 856
rect 114762 2 114870 856
rect 115038 2 115238 856
rect 115406 2 115606 856
rect 115774 2 115974 856
rect 116142 2 116342 856
rect 116510 2 116710 856
rect 116878 2 117078 856
rect 117246 2 117446 856
rect 117614 2 117814 856
rect 117982 2 118182 856
rect 118350 2 118550 856
rect 118718 2 118918 856
rect 119086 2 119286 856
rect 119454 2 119654 856
rect 119822 2 120022 856
rect 120190 2 120390 856
rect 120558 2 120758 856
rect 120926 2 121126 856
rect 121294 2 121494 856
rect 121662 2 121862 856
rect 122030 2 122230 856
rect 122398 2 122598 856
rect 122766 2 122966 856
rect 123134 2 123334 856
rect 123502 2 123702 856
rect 123870 2 124070 856
rect 124238 2 124438 856
rect 124606 2 124806 856
rect 124974 2 125174 856
rect 125342 2 125542 856
rect 125710 2 125910 856
rect 126078 2 126278 856
rect 126446 2 126646 856
rect 126814 2 127014 856
rect 127182 2 127382 856
rect 127550 2 127750 856
rect 127918 2 128118 856
rect 128286 2 128486 856
rect 128654 2 128854 856
rect 129022 2 129222 856
rect 129390 2 129590 856
rect 129758 2 129958 856
rect 130126 2 130326 856
rect 130494 2 130694 856
rect 130862 2 130970 856
rect 131138 2 131338 856
rect 131506 2 131706 856
rect 131874 2 132074 856
rect 132242 2 132442 856
rect 132610 2 132810 856
rect 132978 2 133178 856
rect 133346 2 133546 856
rect 133714 2 133914 856
rect 134082 2 134282 856
rect 134450 2 134650 856
rect 134818 2 135018 856
rect 135186 2 135386 856
rect 135554 2 135754 856
rect 135922 2 136122 856
rect 136290 2 136490 856
rect 136658 2 136858 856
rect 137026 2 137226 856
rect 137394 2 137594 856
rect 137762 2 137962 856
rect 138130 2 138330 856
rect 138498 2 138698 856
rect 138866 2 139066 856
rect 139234 2 139434 856
rect 139602 2 139802 856
rect 139970 2 140170 856
rect 140338 2 140538 856
rect 140706 2 140906 856
rect 141074 2 141274 856
rect 141442 2 141642 856
rect 141810 2 142010 856
rect 142178 2 142378 856
rect 142546 2 142746 856
rect 142914 2 143114 856
rect 143282 2 143482 856
rect 143650 2 143850 856
rect 144018 2 144218 856
rect 144386 2 144586 856
rect 144754 2 144954 856
rect 145122 2 145322 856
rect 145490 2 145690 856
rect 145858 2 146058 856
rect 146226 2 146426 856
rect 146594 2 146794 856
rect 146962 2 147162 856
rect 147330 2 147438 856
rect 147606 2 147806 856
rect 147974 2 148174 856
rect 148342 2 148542 856
rect 148710 2 148910 856
rect 149078 2 149278 856
rect 149446 2 149646 856
rect 149814 2 150014 856
rect 150182 2 150382 856
rect 150550 2 150750 856
rect 150918 2 151118 856
rect 151286 2 151486 856
rect 151654 2 151854 856
rect 152022 2 152222 856
rect 152390 2 152590 856
rect 152758 2 152958 856
rect 153126 2 153326 856
rect 153494 2 153694 856
rect 153862 2 154062 856
rect 154230 2 154430 856
rect 154598 2 154798 856
rect 154966 2 155166 856
rect 155334 2 155534 856
rect 155702 2 155902 856
rect 156070 2 156270 856
rect 156438 2 156638 856
rect 156806 2 157006 856
rect 157174 2 157374 856
rect 157542 2 157742 856
rect 157910 2 158110 856
rect 158278 2 158478 856
rect 158646 2 158846 856
rect 159014 2 159214 856
rect 159382 2 159582 856
rect 159750 2 159950 856
rect 160118 2 160318 856
rect 160486 2 160686 856
rect 160854 2 161054 856
rect 161222 2 161422 856
rect 161590 2 161790 856
rect 161958 2 162158 856
rect 162326 2 162526 856
rect 162694 2 162894 856
rect 163062 2 163262 856
rect 163430 2 163630 856
rect 163798 2 163906 856
rect 164074 2 164274 856
rect 164442 2 164642 856
rect 164810 2 165010 856
rect 165178 2 165378 856
rect 165546 2 165746 856
rect 165914 2 166114 856
rect 166282 2 166482 856
rect 166650 2 166850 856
rect 167018 2 167218 856
rect 167386 2 167586 856
rect 167754 2 167954 856
rect 168122 2 168322 856
rect 168490 2 168690 856
rect 168858 2 169058 856
rect 169226 2 169426 856
rect 169594 2 169794 856
rect 169962 2 170162 856
rect 170330 2 170530 856
rect 170698 2 170898 856
rect 171066 2 171266 856
rect 171434 2 171634 856
rect 171802 2 172002 856
rect 172170 2 172370 856
rect 172538 2 172738 856
rect 172906 2 173106 856
rect 173274 2 173474 856
rect 173642 2 173842 856
rect 174010 2 174210 856
rect 174378 2 174578 856
rect 174746 2 174946 856
rect 175114 2 175314 856
rect 175482 2 175682 856
rect 175850 2 176050 856
rect 176218 2 176418 856
rect 176586 2 176786 856
rect 176954 2 177154 856
rect 177322 2 177522 856
rect 177690 2 177890 856
rect 178058 2 178258 856
rect 178426 2 178626 856
rect 178794 2 178994 856
rect 179162 2 179362 856
rect 179530 2 179730 856
<< obsm3 >>
rect 2221 35 176535 117537
<< metal4 >>
rect 4208 2128 4528 117552
rect 4868 2176 5188 117504
rect 5528 2176 5848 117504
rect 6188 2176 6508 117504
rect 19568 2128 19888 117552
rect 20228 2176 20548 117504
rect 20888 2176 21208 117504
rect 21548 2176 21868 117504
rect 34928 2128 35248 117552
rect 35588 2176 35908 117504
rect 36248 2176 36568 117504
rect 36908 2176 37228 117504
rect 50288 2128 50608 117552
rect 50948 2176 51268 117504
rect 51608 2176 51928 117504
rect 52268 2176 52588 117504
rect 65648 2128 65968 117552
rect 66308 2176 66628 117504
rect 66968 2176 67288 117504
rect 67628 2176 67948 117504
rect 81008 2128 81328 117552
rect 81668 2176 81988 117504
rect 82328 2176 82648 117504
rect 82988 2176 83308 117504
rect 96368 2128 96688 117552
rect 97028 2176 97348 117504
rect 97688 2176 98008 117504
rect 98348 2176 98668 117504
rect 111728 2128 112048 117552
rect 112388 2176 112708 117504
rect 113048 2176 113368 117504
rect 113708 2176 114028 117504
rect 127088 2128 127408 117552
rect 127748 2176 128068 117504
rect 128408 2176 128728 117504
rect 129068 2176 129388 117504
rect 142448 2128 142768 117552
rect 143108 2176 143428 117504
rect 143768 2176 144088 117504
rect 144428 2176 144748 117504
rect 157808 2128 158128 117552
rect 158468 2176 158788 117504
rect 159128 2176 159448 117504
rect 159788 2176 160108 117504
rect 173168 2128 173488 117552
rect 173828 2176 174148 117504
rect 174488 2176 174808 117504
rect 175148 2176 175468 117504
<< obsm4 >>
rect 24998 2048 34848 75309
rect 35328 2096 35508 75309
rect 35988 2096 36168 75309
rect 36648 2096 36828 75309
rect 37308 2096 50208 75309
rect 35328 2048 50208 2096
rect 50688 2096 50868 75309
rect 51348 2096 51528 75309
rect 52008 2096 52188 75309
rect 52668 2096 65568 75309
rect 50688 2048 65568 2096
rect 66048 2096 66228 75309
rect 66708 2096 66888 75309
rect 67368 2096 67548 75309
rect 68028 2096 80928 75309
rect 66048 2048 80928 2096
rect 81408 2096 81588 75309
rect 82068 2096 82248 75309
rect 82728 2096 82908 75309
rect 83388 2096 96288 75309
rect 81408 2048 96288 2096
rect 96768 2096 96948 75309
rect 97428 2096 97608 75309
rect 98088 2096 98268 75309
rect 98748 2096 111648 75309
rect 96768 2048 111648 2096
rect 112128 2096 112308 75309
rect 112788 2096 112968 75309
rect 113448 2096 113628 75309
rect 114108 2096 127008 75309
rect 112128 2048 127008 2096
rect 127488 2096 127668 75309
rect 128148 2096 128328 75309
rect 128808 2096 128988 75309
rect 129468 2096 142368 75309
rect 127488 2048 142368 2096
rect 142848 2096 143028 75309
rect 143508 2096 143688 75309
rect 144168 2096 144348 75309
rect 144828 2096 154317 75309
rect 142848 2048 154317 2096
rect 24998 35 154317 2048
<< obsm5 >>
rect 24956 2900 89860 4580
<< labels >>
rlabel metal2 s 754 119200 810 120000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 47674 119200 47730 120000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 52366 119200 52422 120000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 57058 119200 57114 120000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 61750 119200 61806 120000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 66442 119200 66498 120000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 71134 119200 71190 120000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 75826 119200 75882 120000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 80518 119200 80574 120000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 85210 119200 85266 120000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 89902 119200 89958 120000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 5446 119200 5502 120000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 94686 119200 94742 120000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 99378 119200 99434 120000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 104070 119200 104126 120000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 108762 119200 108818 120000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 113454 119200 113510 120000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 118146 119200 118202 120000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 122838 119200 122894 120000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 127530 119200 127586 120000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 132222 119200 132278 120000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 136914 119200 136970 120000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 10138 119200 10194 120000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 141606 119200 141662 120000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 146298 119200 146354 120000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 150990 119200 151046 120000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 155682 119200 155738 120000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 160374 119200 160430 120000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 165066 119200 165122 120000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 169758 119200 169814 120000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 174450 119200 174506 120000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 14830 119200 14886 120000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 19522 119200 19578 120000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 24214 119200 24270 120000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 28906 119200 28962 120000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 33598 119200 33654 120000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 38290 119200 38346 120000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 42982 119200 43038 120000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 2318 119200 2374 120000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 49238 119200 49294 120000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 53930 119200 53986 120000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 58622 119200 58678 120000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 63314 119200 63370 120000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 68006 119200 68062 120000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 72698 119200 72754 120000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 77390 119200 77446 120000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 82082 119200 82138 120000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 86774 119200 86830 120000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 91558 119200 91614 120000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 7010 119200 7066 120000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 96250 119200 96306 120000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 100942 119200 100998 120000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 105634 119200 105690 120000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 110326 119200 110382 120000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 115018 119200 115074 120000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 119710 119200 119766 120000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 124402 119200 124458 120000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 129094 119200 129150 120000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 133786 119200 133842 120000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 138478 119200 138534 120000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 11702 119200 11758 120000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 143170 119200 143226 120000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 147862 119200 147918 120000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 152554 119200 152610 120000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 157246 119200 157302 120000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 161938 119200 161994 120000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 166630 119200 166686 120000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 171322 119200 171378 120000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 176014 119200 176070 120000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 16394 119200 16450 120000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 21086 119200 21142 120000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 25778 119200 25834 120000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 30470 119200 30526 120000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 35162 119200 35218 120000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 39854 119200 39910 120000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 44546 119200 44602 120000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 3882 119200 3938 120000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 50802 119200 50858 120000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 55494 119200 55550 120000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 60186 119200 60242 120000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 64878 119200 64934 120000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 69570 119200 69626 120000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 74262 119200 74318 120000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 78954 119200 79010 120000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 83646 119200 83702 120000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 88338 119200 88394 120000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 93122 119200 93178 120000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 8574 119200 8630 120000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 97814 119200 97870 120000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 102506 119200 102562 120000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 107198 119200 107254 120000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 111890 119200 111946 120000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 116582 119200 116638 120000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 121274 119200 121330 120000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 125966 119200 126022 120000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 130658 119200 130714 120000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 135350 119200 135406 120000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 140042 119200 140098 120000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 13266 119200 13322 120000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 144734 119200 144790 120000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 149426 119200 149482 120000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 154118 119200 154174 120000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 158810 119200 158866 120000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 163502 119200 163558 120000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 168194 119200 168250 120000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 172886 119200 172942 120000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 177578 119200 177634 120000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 17958 119200 18014 120000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 22650 119200 22706 120000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 27342 119200 27398 120000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 32034 119200 32090 120000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 36726 119200 36782 120000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 41418 119200 41474 120000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 46110 119200 46166 120000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 179418 0 179474 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 179142 119200 179198 120000 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 179786 0 179842 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 38842 0 38898 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 148598 0 148654 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 149702 0 149758 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 150806 0 150862 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 151910 0 151966 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 153014 0 153070 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 154118 0 154174 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 155222 0 155278 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 156326 0 156382 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 157430 0 157486 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 158534 0 158590 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 159638 0 159694 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 160742 0 160798 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 161846 0 161902 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 162950 0 163006 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 163962 0 164018 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 165066 0 165122 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 166170 0 166226 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 167274 0 167330 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 168378 0 168434 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 169482 0 169538 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 170586 0 170642 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 171690 0 171746 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 172794 0 172850 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 173898 0 173954 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 175002 0 175058 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 176106 0 176162 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 177210 0 177266 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 178314 0 178370 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 51998 0 52054 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 54206 0 54262 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 55310 0 55366 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 56414 0 56470 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 57518 0 57574 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 59726 0 59782 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 60830 0 60886 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 61934 0 61990 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 64142 0 64198 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 65246 0 65302 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 66258 0 66314 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 67362 0 67418 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 68466 0 68522 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 70674 0 70730 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 41050 0 41106 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 71778 0 71834 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 72882 0 72938 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 73986 0 74042 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 75090 0 75146 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 76194 0 76250 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 77298 0 77354 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 78402 0 78458 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 79506 0 79562 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 80610 0 80666 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 81714 0 81770 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 42154 0 42210 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 82726 0 82782 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 83830 0 83886 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 84934 0 84990 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 86038 0 86094 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 87142 0 87198 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 89350 0 89406 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 90454 0 90510 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 92662 0 92718 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 93766 0 93822 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 95974 0 96030 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 98182 0 98238 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 99194 0 99250 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 100298 0 100354 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 101402 0 101458 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 102506 0 102562 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 103610 0 103666 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 44362 0 44418 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 104714 0 104770 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 105818 0 105874 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 106922 0 106978 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 108026 0 108082 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 109130 0 109186 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 110234 0 110290 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 111338 0 111394 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 112442 0 112498 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 113546 0 113602 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 114650 0 114706 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 115662 0 115718 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 116766 0 116822 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 117870 0 117926 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 118974 0 119030 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 120078 0 120134 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 121182 0 121238 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 122286 0 122342 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 123390 0 123446 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 124494 0 124550 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 125598 0 125654 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 126702 0 126758 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 127806 0 127862 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 128910 0 128966 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 130014 0 130070 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 131026 0 131082 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 132130 0 132186 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 133234 0 133290 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 134338 0 134394 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 135442 0 135498 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 136546 0 136602 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 137650 0 137706 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 138754 0 138810 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 139858 0 139914 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 140962 0 141018 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 142066 0 142122 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 143170 0 143226 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 144274 0 144330 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 145378 0 145434 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 146482 0 146538 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 147494 0 147550 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 48778 0 48834 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 148966 0 149022 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 150070 0 150126 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 151174 0 151230 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 152278 0 152334 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 153382 0 153438 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 154486 0 154542 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 155590 0 155646 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 156694 0 156750 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 157798 0 157854 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 158902 0 158958 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 50158 0 50214 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 160006 0 160062 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 161110 0 161166 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 162214 0 162270 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 163318 0 163374 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 164330 0 164386 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 165434 0 165490 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 166538 0 166594 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 167642 0 167698 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 168746 0 168802 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 169850 0 169906 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 51262 0 51318 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 170954 0 171010 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 172058 0 172114 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 173162 0 173218 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 174266 0 174322 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 175370 0 175426 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 176474 0 176530 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 177578 0 177634 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 178682 0 178738 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 52366 0 52422 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 53470 0 53526 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 54574 0 54630 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 55678 0 55734 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 56782 0 56838 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 57886 0 57942 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 58990 0 59046 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 60094 0 60150 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 40314 0 40370 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 61198 0 61254 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 62302 0 62358 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 63406 0 63462 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 64510 0 64566 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 65522 0 65578 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 66626 0 66682 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 67730 0 67786 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 68834 0 68890 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 69938 0 69994 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 71042 0 71098 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 41418 0 41474 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 72146 0 72202 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 73250 0 73306 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 74354 0 74410 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 75458 0 75514 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 76562 0 76618 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 77666 0 77722 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 78770 0 78826 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 79874 0 79930 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 80978 0 81034 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 81990 0 82046 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 42522 0 42578 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 83094 0 83150 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 84198 0 84254 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 85302 0 85358 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 86406 0 86462 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 87510 0 87566 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 88614 0 88670 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 89718 0 89774 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 90822 0 90878 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 91926 0 91982 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 93030 0 93086 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 43626 0 43682 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 94134 0 94190 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 95238 0 95294 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 96342 0 96398 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 97446 0 97502 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 98458 0 98514 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 99562 0 99618 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 100666 0 100722 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 101770 0 101826 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 102874 0 102930 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 103978 0 104034 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 44730 0 44786 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 105082 0 105138 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 106186 0 106242 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 107290 0 107346 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 108394 0 108450 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 109498 0 109554 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 110602 0 110658 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 111706 0 111762 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 112810 0 112866 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 113914 0 113970 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 114926 0 114982 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 45834 0 45890 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 116030 0 116086 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 117134 0 117190 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 118238 0 118294 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 119342 0 119398 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 120446 0 120502 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 121550 0 121606 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 122654 0 122710 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 123758 0 123814 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 124862 0 124918 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 125966 0 126022 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 46938 0 46994 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 127070 0 127126 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 128174 0 128230 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 129278 0 129334 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 130382 0 130438 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 131394 0 131450 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 132498 0 132554 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 133602 0 133658 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 134706 0 134762 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 135810 0 135866 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 136914 0 136970 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 48042 0 48098 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 138018 0 138074 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 139122 0 139178 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 140226 0 140282 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 141330 0 141386 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 142434 0 142490 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 143538 0 143594 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 144642 0 144698 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 145746 0 145802 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 146850 0 146906 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 147862 0 147918 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 49146 0 49202 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 39578 0 39634 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 149334 0 149390 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 150438 0 150494 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 151542 0 151598 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 152646 0 152702 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 153750 0 153806 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 154854 0 154910 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 155958 0 156014 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 157062 0 157118 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 158166 0 158222 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 159270 0 159326 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 50526 0 50582 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 160374 0 160430 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 161478 0 161534 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 162582 0 162638 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 163686 0 163742 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 164698 0 164754 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 165802 0 165858 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 166906 0 166962 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 168010 0 168066 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 169114 0 169170 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 170218 0 170274 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 51630 0 51686 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 171322 0 171378 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 172426 0 172482 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 173530 0 173586 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 174634 0 174690 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 175738 0 175794 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 176842 0 176898 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 177946 0 178002 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 179050 0 179106 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 57150 0 57206 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 58254 0 58310 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 40682 0 40738 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 61566 0 61622 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 62670 0 62726 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 64878 0 64934 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 65890 0 65946 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 68098 0 68154 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 69202 0 69258 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 70306 0 70362 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 71410 0 71466 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 41786 0 41842 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 72514 0 72570 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 73618 0 73674 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 74722 0 74778 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 75826 0 75882 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 78034 0 78090 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 80242 0 80298 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 81346 0 81402 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 83462 0 83518 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 84566 0 84622 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 85670 0 85726 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 86774 0 86830 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 88982 0 89038 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 90086 0 90142 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 91190 0 91246 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 92294 0 92350 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 43994 0 44050 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 94502 0 94558 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 95606 0 95662 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 96710 0 96766 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 97814 0 97870 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 98826 0 98882 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 99930 0 99986 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 101034 0 101090 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 102138 0 102194 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 103242 0 103298 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 104346 0 104402 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 105450 0 105506 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 106554 0 106610 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 107658 0 107714 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 108762 0 108818 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 109866 0 109922 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 110970 0 111026 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 112074 0 112130 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 113178 0 113234 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 114282 0 114338 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 115294 0 115350 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 46202 0 46258 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 116398 0 116454 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 117502 0 117558 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 118606 0 118662 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 119710 0 119766 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 120814 0 120870 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 121918 0 121974 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 123022 0 123078 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 124126 0 124182 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 125230 0 125286 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 126334 0 126390 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 127438 0 127494 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 128542 0 128598 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 129646 0 129702 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 130750 0 130806 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 131762 0 131818 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 132866 0 132922 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 133970 0 134026 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 135074 0 135130 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 136178 0 136234 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 137282 0 137338 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 48410 0 48466 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 138386 0 138442 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 139490 0 139546 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 140594 0 140650 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 141698 0 141754 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 142802 0 142858 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 143906 0 143962 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 145010 0 145066 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 146114 0 146170 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 147218 0 147274 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 148230 0 148286 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 502 nsew signal input
rlabel metal2 s 386 0 442 800 6 wb_rst_i
port 503 nsew signal input
rlabel metal2 s 754 0 810 800 6 wbs_ack_o
port 504 nsew signal output
rlabel metal2 s 2226 0 2282 800 6 wbs_adr_i[0]
port 505 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 wbs_adr_i[10]
port 506 nsew signal input
rlabel metal2 s 15842 0 15898 800 6 wbs_adr_i[11]
port 507 nsew signal input
rlabel metal2 s 16854 0 16910 800 6 wbs_adr_i[12]
port 508 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 wbs_adr_i[13]
port 509 nsew signal input
rlabel metal2 s 19062 0 19118 800 6 wbs_adr_i[14]
port 510 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 wbs_adr_i[15]
port 511 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 wbs_adr_i[16]
port 512 nsew signal input
rlabel metal2 s 22374 0 22430 800 6 wbs_adr_i[17]
port 513 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 wbs_adr_i[18]
port 514 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 wbs_adr_i[19]
port 515 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_adr_i[1]
port 516 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 wbs_adr_i[20]
port 517 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 wbs_adr_i[21]
port 518 nsew signal input
rlabel metal2 s 27894 0 27950 800 6 wbs_adr_i[22]
port 519 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 wbs_adr_i[23]
port 520 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 wbs_adr_i[24]
port 521 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 wbs_adr_i[25]
port 522 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 wbs_adr_i[26]
port 523 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 wbs_adr_i[27]
port 524 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 wbs_adr_i[28]
port 525 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 wbs_adr_i[29]
port 526 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_adr_i[2]
port 527 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 wbs_adr_i[30]
port 528 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 wbs_adr_i[31]
port 529 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 wbs_adr_i[3]
port 530 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_adr_i[4]
port 531 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 wbs_adr_i[5]
port 532 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wbs_adr_i[6]
port 533 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 wbs_adr_i[7]
port 534 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 wbs_adr_i[8]
port 535 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 wbs_adr_i[9]
port 536 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wbs_cyc_i
port 537 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_dat_i[0]
port 538 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 wbs_dat_i[10]
port 539 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 wbs_dat_i[11]
port 540 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 wbs_dat_i[12]
port 541 nsew signal input
rlabel metal2 s 18326 0 18382 800 6 wbs_dat_i[13]
port 542 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 wbs_dat_i[14]
port 543 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 wbs_dat_i[15]
port 544 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 wbs_dat_i[16]
port 545 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 wbs_dat_i[17]
port 546 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 wbs_dat_i[18]
port 547 nsew signal input
rlabel metal2 s 24950 0 25006 800 6 wbs_dat_i[19]
port 548 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 wbs_dat_i[1]
port 549 nsew signal input
rlabel metal2 s 26054 0 26110 800 6 wbs_dat_i[20]
port 550 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 wbs_dat_i[21]
port 551 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 wbs_dat_i[22]
port 552 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 wbs_dat_i[23]
port 553 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 wbs_dat_i[24]
port 554 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 wbs_dat_i[25]
port 555 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 wbs_dat_i[26]
port 556 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 wbs_dat_i[27]
port 557 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 wbs_dat_i[28]
port 558 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 wbs_dat_i[29]
port 559 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 wbs_dat_i[2]
port 560 nsew signal input
rlabel metal2 s 37002 0 37058 800 6 wbs_dat_i[30]
port 561 nsew signal input
rlabel metal2 s 38106 0 38162 800 6 wbs_dat_i[31]
port 562 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 wbs_dat_i[3]
port 563 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_dat_i[4]
port 564 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_i[5]
port 565 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 wbs_dat_i[6]
port 566 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 wbs_dat_i[7]
port 567 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 wbs_dat_i[8]
port 568 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 wbs_dat_i[9]
port 569 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 wbs_dat_o[0]
port 570 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 wbs_dat_o[10]
port 571 nsew signal output
rlabel metal2 s 16486 0 16542 800 6 wbs_dat_o[11]
port 572 nsew signal output
rlabel metal2 s 17590 0 17646 800 6 wbs_dat_o[12]
port 573 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 wbs_dat_o[13]
port 574 nsew signal output
rlabel metal2 s 19798 0 19854 800 6 wbs_dat_o[14]
port 575 nsew signal output
rlabel metal2 s 20902 0 20958 800 6 wbs_dat_o[15]
port 576 nsew signal output
rlabel metal2 s 22006 0 22062 800 6 wbs_dat_o[16]
port 577 nsew signal output
rlabel metal2 s 23110 0 23166 800 6 wbs_dat_o[17]
port 578 nsew signal output
rlabel metal2 s 24214 0 24270 800 6 wbs_dat_o[18]
port 579 nsew signal output
rlabel metal2 s 25318 0 25374 800 6 wbs_dat_o[19]
port 580 nsew signal output
rlabel metal2 s 4434 0 4490 800 6 wbs_dat_o[1]
port 581 nsew signal output
rlabel metal2 s 26422 0 26478 800 6 wbs_dat_o[20]
port 582 nsew signal output
rlabel metal2 s 27526 0 27582 800 6 wbs_dat_o[21]
port 583 nsew signal output
rlabel metal2 s 28630 0 28686 800 6 wbs_dat_o[22]
port 584 nsew signal output
rlabel metal2 s 29734 0 29790 800 6 wbs_dat_o[23]
port 585 nsew signal output
rlabel metal2 s 30838 0 30894 800 6 wbs_dat_o[24]
port 586 nsew signal output
rlabel metal2 s 31942 0 31998 800 6 wbs_dat_o[25]
port 587 nsew signal output
rlabel metal2 s 32954 0 33010 800 6 wbs_dat_o[26]
port 588 nsew signal output
rlabel metal2 s 34058 0 34114 800 6 wbs_dat_o[27]
port 589 nsew signal output
rlabel metal2 s 35162 0 35218 800 6 wbs_dat_o[28]
port 590 nsew signal output
rlabel metal2 s 36266 0 36322 800 6 wbs_dat_o[29]
port 591 nsew signal output
rlabel metal2 s 5906 0 5962 800 6 wbs_dat_o[2]
port 592 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 wbs_dat_o[30]
port 593 nsew signal output
rlabel metal2 s 38474 0 38530 800 6 wbs_dat_o[31]
port 594 nsew signal output
rlabel metal2 s 7378 0 7434 800 6 wbs_dat_o[3]
port 595 nsew signal output
rlabel metal2 s 8850 0 8906 800 6 wbs_dat_o[4]
port 596 nsew signal output
rlabel metal2 s 9954 0 10010 800 6 wbs_dat_o[5]
port 597 nsew signal output
rlabel metal2 s 11058 0 11114 800 6 wbs_dat_o[6]
port 598 nsew signal output
rlabel metal2 s 12162 0 12218 800 6 wbs_dat_o[7]
port 599 nsew signal output
rlabel metal2 s 13266 0 13322 800 6 wbs_dat_o[8]
port 600 nsew signal output
rlabel metal2 s 14370 0 14426 800 6 wbs_dat_o[9]
port 601 nsew signal output
rlabel metal2 s 3330 0 3386 800 6 wbs_sel_i[0]
port 602 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 wbs_sel_i[1]
port 603 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 wbs_sel_i[2]
port 604 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wbs_sel_i[3]
port 605 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_stb_i
port 606 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 wbs_we_i
port 607 nsew signal input
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 608 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 609 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 610 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 611 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 612 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 613 nsew power bidirectional
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 614 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 615 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 616 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 617 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 618 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 619 nsew ground bidirectional
rlabel metal4 s 158468 2176 158788 117504 6 vccd2
port 620 nsew power bidirectional
rlabel metal4 s 127748 2176 128068 117504 6 vccd2
port 621 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 117504 6 vccd2
port 622 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 117504 6 vccd2
port 623 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 117504 6 vccd2
port 624 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 117504 6 vccd2
port 625 nsew power bidirectional
rlabel metal4 s 173828 2176 174148 117504 6 vssd2
port 626 nsew ground bidirectional
rlabel metal4 s 143108 2176 143428 117504 6 vssd2
port 627 nsew ground bidirectional
rlabel metal4 s 112388 2176 112708 117504 6 vssd2
port 628 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 117504 6 vssd2
port 629 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 117504 6 vssd2
port 630 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 117504 6 vssd2
port 631 nsew ground bidirectional
rlabel metal4 s 159128 2176 159448 117504 6 vdda1
port 632 nsew power bidirectional
rlabel metal4 s 128408 2176 128728 117504 6 vdda1
port 633 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 117504 6 vdda1
port 634 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 117504 6 vdda1
port 635 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 117504 6 vdda1
port 636 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 117504 6 vdda1
port 637 nsew power bidirectional
rlabel metal4 s 174488 2176 174808 117504 6 vssa1
port 638 nsew ground bidirectional
rlabel metal4 s 143768 2176 144088 117504 6 vssa1
port 639 nsew ground bidirectional
rlabel metal4 s 113048 2176 113368 117504 6 vssa1
port 640 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 117504 6 vssa1
port 641 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 117504 6 vssa1
port 642 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 117504 6 vssa1
port 643 nsew ground bidirectional
rlabel metal4 s 159788 2176 160108 117504 6 vdda2
port 644 nsew power bidirectional
rlabel metal4 s 129068 2176 129388 117504 6 vdda2
port 645 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 117504 6 vdda2
port 646 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 117504 6 vdda2
port 647 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 117504 6 vdda2
port 648 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 117504 6 vdda2
port 649 nsew power bidirectional
rlabel metal4 s 175148 2176 175468 117504 6 vssa2
port 650 nsew ground bidirectional
rlabel metal4 s 144428 2176 144748 117504 6 vssa2
port 651 nsew ground bidirectional
rlabel metal4 s 113708 2176 114028 117504 6 vssa2
port 652 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 117504 6 vssa2
port 653 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 117504 6 vssa2
port 654 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 117504 6 vssa2
port 655 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 180000 120000
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
string GDS_END 51412460
string GDS_START 1373928
<< end >>

